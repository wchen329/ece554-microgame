module audio_controller(
	input clk, rst_n,
	input set_tone,
	input [31:0] tone
);

endmodule
