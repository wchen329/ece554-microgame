// soc_audio.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_audio (
		input  wire [1:0]  address,     // avalon_audio_slave.address
		input  wire        chipselect,  //                   .chipselect
		input  wire        read,        //                   .read
		input  wire        write,       //                   .write
		input  wire [31:0] writedata,   //                   .writedata
		output wire [31:0] readdata,    //                   .readdata
		input  wire        clk,         //                clk.clk
		input  wire        AUD_BCLK,    // external_interface.BCLK
		output wire        AUD_DACDAT,  //                   .DACDAT
		input  wire        AUD_DACLRCK, //                   .DACLRCK
		output wire        irq,         //          interrupt.irq
		input  wire        reset        //              reset.reset
	);

	soc_audio_audio_0 audio_0 (
		.clk         (clk),         //                clk.clk
		.reset       (reset),       //              reset.reset
		.address     (address),     // avalon_audio_slave.address
		.chipselect  (chipselect),  //                   .chipselect
		.read        (read),        //                   .read
		.write       (write),       //                   .write
		.writedata   (writedata),   //                   .writedata
		.readdata    (readdata),    //                   .readdata
		.irq         (irq),         //          interrupt.irq
		.AUD_BCLK    (AUD_BCLK),    // external_interface.export
		.AUD_DACDAT  (AUD_DACDAT),  //                   .export
		.AUD_DACLRCK (AUD_DACLRCK)  //                   .export
	);

endmodule
