module input_buffer(
	input clk, rst_n,
	input clear,
	input up, right, down, left, space
);

endmodule
