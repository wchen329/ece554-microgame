
// logic [27:0] stim_mem [1000];
// $readmemh("files/band_scale_stim.hex", stim_mem);