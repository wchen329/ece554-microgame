module sprite_command_fifo_front_end(
	input clk, rst_n,
	input [79:0] cmd,
	input write
);

endmodule
