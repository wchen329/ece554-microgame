module instruction_memory
#(
	parameter DATA_WIDTH_BLAH_BLAH_BLAH=16,
	localparam MAX_INSTRUCTIONS=256
)(
	input clk,
	input [15:0] address_a, address_b,
	output [31:0] data_a, data_b
);

int fd;

integer i;
reg [31:0] instructions[MAX_INSTRUCTIONS-1:0];

reg [31:0] addr;

always_ff @(posedge clk) begin
	addr <= {21'b0, address_a[10:0]};
end


// read in fake instuction memory file
// make sure to add delay so this can complete
initial begin
	fd = $fopen("ece554-microgame/v/testing/cpu_test_harness/instructions.hl", "r");

	if(fd == 0) begin
		$display("Could not open file");
		$finish();
	end

	// clear memory
	for(i=0; i<MAX_INSTRUCTIONS; i=i+1) begin
		instructions[i] = 32'b0;
	end

	i = 0;
	while(i<MAX_INSTRUCTIONS && ~$feof(fd) && $fscanf(fd, "%h\n", instructions[i]) == 1) begin
		$display("loaded instruction: %b", instructions[i]);
		i = i + 1;
	end

	$fclose(fd);
end

assign data_a = addr >= MAX_INSTRUCTIONS ? 32'b0 : instructions[addr];

assign data_b = 16'h0000;

endmodule
