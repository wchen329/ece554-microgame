LOOP:
lk $4
b LOOP
