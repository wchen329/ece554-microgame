
module soc_audio_lrclk (
	clk,
	reset,
	AUD_BCLK,
	AUD_LRCLK);	

	input		clk;
	input		reset;
	input		AUD_BCLK;
	output		AUD_LRCLK;
endmodule
